`ifndef CONFIGURATION_PKG_SV
    `define CONFIGURATION_PKG_SV

    package configuration_pkg;

        
        import uvm_pkg::*;     
        `include "uvm_macros.svh" 
        `include "seg_config.sv" 

    endpackage : configuration_pkg

`endif     